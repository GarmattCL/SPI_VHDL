module led (
    input btn1,          // Eingangs-Taster
    output led       // Ausgang-LED
);
assign led = btn1;
endmodule